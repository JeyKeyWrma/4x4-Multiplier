module and_4(A3,A2,A1,A0,B,O3,O2,O1,O0);
    input A3,A2,A1,A0,B;
    output O3,O2,O1,O0;
    and(O3,A3,B);
    and(O2,A2,B);
    and(O1,A1,B);
    and(O0,A0,B);
endmodule

module halfadder(a,b,s,c);

    input a,b;
    output s,c;
    xor sum(s,a,b);
    and carry(c,a,b);
    
endmodule

module fulladder(a,b,c_in,s,c);

    input a,b,c_in;
    output s,c;
    wire n1,n2,n3;

    halfadder adder1(.a(a),.b(b),.s(n1),.c(n2));
    halfadder adder2(.a(c_in),.b(n1),.s(s),.c(n3));
    or carry(c,n2,n3);
    
endmodule

module adder(A3,A2,A1,A0,B3,B2,B1,B0,S4,S3,S2,S1,S0);

    input A3,A2,A1,A0,B3,B2,B1,B0;
    output S4,S3,S2,S1,S0;
    wire n1,n2,n3;
    
    halfadder HA1(A0,B0,S0,n1);
    fulladder FA1(A1,B1,n1,S1,n2);
    fulladder FA2(A2,B2,n2,S2,n3);
    fulladder FA3(A3,B3,n3,S3,S4);
    
endmodule

module multiplier(A3,A2,A1,A0,B3,B2,B1,B0,p7,p6,p5,p4,p3,p2,p1,p0);

    input A3,A2,A1,A0,B3,B2,B1,B0;
    output p7,p6,p5,p4,p3,p2,p1,p0;
    wire n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,n20,n21,n22,n23,temp; 

    assign temp =0;
    and_4 AL1(A3,A2,A1,A0,B0,n1,n2,n3,p0);

    and_4 AL2(A3,A2,A1,A0,B1,n4,n5,n6,n7);
    adder ad1(temp,n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,p1);

    and_4 AL3(A3,A2,A1,A0,B2,n12,n13,n14,n15);
    adder ad2(n8,n9,n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,p2);

    and_4 AL4(A3,A2,A1,A0,B3,n20,n21,n22,n23);
    adder ad3(n16,n17,n18,n19,n20,n21,n22,n23,p7,p6,p5,p4,p3);


endmodule

module testbench;
wire [7:0]P;
reg [3:0] A,B;

multiplier my_gate(A[3],A[2],A[1],A[0],B[3],B[2],B[1],B[0],P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0]);

initial
begin
    $dumpfile("runfile.vcd");
    $dumpvars(0,testbench);
    A = 4'b0000;
    B = 4'b0000;
end
initial 
begin
$monitor("inputs A= ",A,"\ninputs B= ",B,"\noutput = ",P[7],P[6],P[5],P[4],P[3],P[2],P[1],P[0]);

A = 4'b0000;
B = 4'b0000;
#5
A = 4'b0000;
B = 4'b0001;
#5
A = 4'b0000;
B = 4'b0010;
#5
A = 4'b0000;
B = 4'b0011;
#5
A = 4'b0000;
B = 4'b0100;
#5
A = 4'b0000;
B = 4'b0101;
#5
A = 4'b0000;
B = 4'b0110;
#5
A = 4'b0000;
B = 4'b0111;
#5
A = 4'b0000;
B = 4'b1000;
#5
A = 4'b0000;
B = 4'b1001;
#5
A = 4'b0000;
B = 4'b1010;
#5
A = 4'b0000;
B = 4'b1011;
#5
A = 4'b0000;
B = 4'b1100;
#5
A = 4'b0000;
B = 4'b1101;
#5
A = 4'b0000;
B = 4'b1110;
#5
A = 4'b0000;
B = 4'b1111;
#5
A = 4'b0001;
B = 4'b0000;
#5
A = 4'b0001;
B = 4'b0001;
#5
A = 4'b0001;
B = 4'b0010;
#5
A = 4'b0001;
B = 4'b0011;
#5
A = 4'b0001;
B = 4'b0100;
#5
A = 4'b0001;
B = 4'b0101;
#5
A = 4'b0001;
B = 4'b0110;
#5
A = 4'b0001;
B = 4'b0111;
#5
A = 4'b0001;
B = 4'b1000;
#5
A = 4'b0001;
B = 4'b1001;
#5
A = 4'b0001;
B = 4'b1010;
#5
A = 4'b0001;
B = 4'b1011;
#5
A = 4'b0001;
B = 4'b1100;
#5
A = 4'b0001;
B = 4'b1101;
#5
A = 4'b0001;
B = 4'b1110;
#5
A = 4'b0001;
B = 4'b1111;
#5
A = 4'b0010;
B = 4'b0000;
#5
A = 4'b0010;
B = 4'b0001;
#5
A = 4'b0010;
B = 4'b0010;
#5
A = 4'b0010;
B = 4'b0011;
#5
A = 4'b0010;
B = 4'b0100;
#5
A = 4'b0010;
B = 4'b0101;
#5
A = 4'b0010;
B = 4'b0110;
#5
A = 4'b0010;
B = 4'b0111;
#5
A = 4'b0010;
B = 4'b1000;
#5
A = 4'b0010;
B = 4'b1001;
#5
A = 4'b0010;
B = 4'b1010;
#5
A = 4'b0010;
B = 4'b1011;
#5
A = 4'b0010;
B = 4'b1100;
#5
A = 4'b0010;
B = 4'b1101;
#5
A = 4'b0010;
B = 4'b1110;
#5
A = 4'b0010;
B = 4'b1111;
#5
A = 4'b0011;
B = 4'b0000;
#5
A = 4'b0011;
B = 4'b0001;
#5
A = 4'b0011;
B = 4'b0010;
#5
A = 4'b0011;
B = 4'b0011;
#5
A = 4'b0011;
B = 4'b0100;
#5
A = 4'b0011;
B = 4'b0101;
#5
A = 4'b0011;
B = 4'b0110;
#5
A = 4'b0011;
B = 4'b0111;
#5
A = 4'b0011;
B = 4'b1000;
#5
A = 4'b0011;
B = 4'b1001;
#5
A = 4'b0011;
B = 4'b1010;
#5
A = 4'b0011;
B = 4'b1011;
#5
A = 4'b0011;
B = 4'b1100;
#5
A = 4'b0011;
B = 4'b1101;
#5
A = 4'b0011;
B = 4'b1110;
#5
A = 4'b0011;
B = 4'b1111;
#5
A = 4'b0100;
B = 4'b0000;
#5
A = 4'b0100;
B = 4'b0001;
#5
A = 4'b0100;
B = 4'b0010;
#5
A = 4'b0100;
B = 4'b0011;
#5
A = 4'b0100;
B = 4'b0100;
#5
A = 4'b0100;
B = 4'b0101;
#5
A = 4'b0100;
B = 4'b0110;
#5
A = 4'b0100;
B = 4'b0111;
#5
A = 4'b0100;
B = 4'b1000;
#5
A = 4'b0100;
B = 4'b1001;
#5
A = 4'b0100;
B = 4'b1010;
#5
A = 4'b0100;
B = 4'b1011;
#5
A = 4'b0100;
B = 4'b1100;
#5
A = 4'b0100;
B = 4'b1101;
#5
A = 4'b0100;
B = 4'b1110;
#5
A = 4'b0100;
B = 4'b1111;
#5
A = 4'b0101;
B = 4'b0000;
#5
A = 4'b0101;
B = 4'b0001;
#5
A = 4'b0101;
B = 4'b0010;
#5
A = 4'b0101;
B = 4'b0011;
#5
A = 4'b0101;
B = 4'b0100;
#5
A = 4'b0101;
B = 4'b0101;
#5
A = 4'b0101;
B = 4'b0110;
#5
A = 4'b0101;
B = 4'b0111;
#5
A = 4'b0101;
B = 4'b1000;
#5
A = 4'b0101;
B = 4'b1001;
#5
A = 4'b0101;
B = 4'b1010;
#5
A = 4'b0101;
B = 4'b1011;
#5
A = 4'b0101;
B = 4'b1100;
#5
A = 4'b0101;
B = 4'b1101;
#5
A = 4'b0101;
B = 4'b1110;
#5
A = 4'b0101;
B = 4'b1111;
#5
A = 4'b0110;
B = 4'b0000;
#5
A = 4'b0110;
B = 4'b0001;
#5
A = 4'b0110;
B = 4'b0010;
#5
A = 4'b0110;
B = 4'b0011;
#5
A = 4'b0110;
B = 4'b0100;
#5
A = 4'b0110;
B = 4'b0101;
#5
A = 4'b0110;
B = 4'b0110;
#5
A = 4'b0110;
B = 4'b0111;
#5
A = 4'b0110;
B = 4'b1000;
#5
A = 4'b0110;
B = 4'b1001;
#5
A = 4'b0110;
B = 4'b1010;
#5
A = 4'b0110;
B = 4'b1011;
#5
A = 4'b0110;
B = 4'b1100;
#5
A = 4'b0110;
B = 4'b1101;
#5
A = 4'b0110;
B = 4'b1110;
#5
A = 4'b0110;
B = 4'b1111;
#5
A = 4'b0111;
B = 4'b0000;
#5
A = 4'b0111;
B = 4'b0001;
#5
A = 4'b0111;
B = 4'b0010;
#5
A = 4'b0111;
B = 4'b0011;
#5
A = 4'b0111;
B = 4'b0100;
#5
A = 4'b0111;
B = 4'b0101;
#5
A = 4'b0111;
B = 4'b0110;
#5
A = 4'b0111;
B = 4'b0111;
#5
A = 4'b0111;
B = 4'b1000;
#5
A = 4'b0111;
B = 4'b1001;
#5
A = 4'b0111;
B = 4'b1010;
#5
A = 4'b0111;
B = 4'b1011;
#5
A = 4'b0111;
B = 4'b1100;
#5
A = 4'b0111;
B = 4'b1101;
#5
A = 4'b0111;
B = 4'b1110;
#5
A = 4'b0111;
B = 4'b1111;
#5
A = 4'b1000;
B = 4'b0000;
#5
A = 4'b1000;
B = 4'b0001;
#5
A = 4'b1000;
B = 4'b0010;
#5
A = 4'b1000;
B = 4'b0011;
#5
A = 4'b1000;
B = 4'b0100;
#5
A = 4'b1000;
B = 4'b0101;
#5
A = 4'b1000;
B = 4'b0110;
#5
A = 4'b1000;
B = 4'b0111;
#5
A = 4'b1000;
B = 4'b1000;
#5
A = 4'b1000;
B = 4'b1001;
#5
A = 4'b1000;
B = 4'b1010;
#5
A = 4'b1000;
B = 4'b1011;
#5
A = 4'b1000;
B = 4'b1100;
#5
A = 4'b1000;
B = 4'b1101;
#5
A = 4'b1000;
B = 4'b1110;
#5
A = 4'b1000;
B = 4'b1111;
#5
A = 4'b1001;
B = 4'b0000;
#5
A = 4'b1001;
B = 4'b0001;
#5
A = 4'b1001;
B = 4'b0010;
#5
A = 4'b1001;
B = 4'b0011;
#5
A = 4'b1001;
B = 4'b0100;
#5
A = 4'b1001;
B = 4'b0101;
#5
A = 4'b1001;
B = 4'b0110;
#5
A = 4'b1001;
B = 4'b0111;
#5
A = 4'b1001;
B = 4'b1000;
#5
A = 4'b1001;
B = 4'b1001;
#5
A = 4'b1001;
B = 4'b1010;
#5
A = 4'b1001;
B = 4'b1011;
#5
A = 4'b1001;
B = 4'b1100;
#5
A = 4'b1001;
B = 4'b1101;
#5
A = 4'b1001;
B = 4'b1110;
#5
A = 4'b1001;
B = 4'b1111;
#5
A = 4'b1010;
B = 4'b0000;
#5
A = 4'b1010;
B = 4'b0001;
#5
A = 4'b1010;
B = 4'b0010;
#5
A = 4'b1010;
B = 4'b0011;
#5
A = 4'b1010;
B = 4'b0100;
#5
A = 4'b1010;
B = 4'b0101;
#5
A = 4'b1010;
B = 4'b0110;
#5
A = 4'b1010;
B = 4'b0111;
#5
A = 4'b1010;
B = 4'b1000;
#5
A = 4'b1010;
B = 4'b1001;
#5
A = 4'b1010;
B = 4'b1010;
#5
A = 4'b1010;
B = 4'b1011;
#5
A = 4'b1010;
B = 4'b1100;
#5
A = 4'b1010;
B = 4'b1101;
#5
A = 4'b1010;
B = 4'b1110;
#5
A = 4'b1010;
B = 4'b1111;
#5
A = 4'b1011;
B = 4'b0000;
#5
A = 4'b1011;
B = 4'b0001;
#5
A = 4'b1011;
B = 4'b0010;
#5
A = 4'b1011;
B = 4'b0011;
#5
A = 4'b1011;
B = 4'b0100;
#5
A = 4'b1011;
B = 4'b0101;
#5
A = 4'b1011;
B = 4'b0110;
#5
A = 4'b1011;
B = 4'b0111;
#5
A = 4'b1011;
B = 4'b1000;
#5
A = 4'b1011;
B = 4'b1001;
#5
A = 4'b1011;
B = 4'b1010;
#5
A = 4'b1011;
B = 4'b1011;
#5
A = 4'b1011;
B = 4'b1100;
#5
A = 4'b1011;
B = 4'b1101;
#5
A = 4'b1011;
B = 4'b1110;
#5
A = 4'b1011;
B = 4'b1111;
#5
A = 4'b1100;
B = 4'b0000;
#5
A = 4'b1100;
B = 4'b0001;
#5
A = 4'b1100;
B = 4'b0010;
#5
A = 4'b1100;
B = 4'b0011;
#5
A = 4'b1100;
B = 4'b0100;
#5
A = 4'b1100;
B = 4'b0101;
#5
A = 4'b1100;
B = 4'b0110;
#5
A = 4'b1100;
B = 4'b0111;
#5
A = 4'b1100;
B = 4'b1000;
#5
A = 4'b1100;
B = 4'b1001;
#5
A = 4'b1100;
B = 4'b1010;
#5
A = 4'b1100;
B = 4'b1011;
#5
A = 4'b1100;
B = 4'b1100;
#5
A = 4'b1100;
B = 4'b1101;
#5
A = 4'b1100;
B = 4'b1110;
#5
A = 4'b1100;
B = 4'b1111;
#5
A = 4'b1101;
B = 4'b0000;
#5
A = 4'b1101;
B = 4'b0001;
#5
A = 4'b1101;
B = 4'b0010;
#5
A = 4'b1101;
B = 4'b0011;
#5
A = 4'b1101;
B = 4'b0100;
#5
A = 4'b1101;
B = 4'b0101;
#5
A = 4'b1101;
B = 4'b0110;
#5
A = 4'b1101;
B = 4'b0111;
#5
A = 4'b1101;
B = 4'b1000;
#5
A = 4'b1101;
B = 4'b1001;
#5
A = 4'b1101;
B = 4'b1010;
#5
A = 4'b1101;
B = 4'b1011;
#5
A = 4'b1101;
B = 4'b1100;
#5
A = 4'b1101;
B = 4'b1101;
#5
A = 4'b1101;
B = 4'b1110;
#5
A = 4'b1101;
B = 4'b1111;
#5
A = 4'b1110;
B = 4'b0000;
#5
A = 4'b1110;
B = 4'b0001;
#5
A = 4'b1110;
B = 4'b0010;
#5
A = 4'b1110;
B = 4'b0011;
#5
A = 4'b1110;
B = 4'b0100;
#5
A = 4'b1110;
B = 4'b0101;
#5
A = 4'b1110;
B = 4'b0110;
#5
A = 4'b1110;
B = 4'b0111;
#5
A = 4'b1110;
B = 4'b1000;
#5
A = 4'b1110;
B = 4'b1001;
#5
A = 4'b1110;
B = 4'b1010;
#5
A = 4'b1110;
B = 4'b1011;
#5
A = 4'b1110;
B = 4'b1100;
#5
A = 4'b1110;
B = 4'b1101;
#5
A = 4'b1110;
B = 4'b1110;
#5
A = 4'b1110;
B = 4'b1111;
#5
A = 4'b1111;
B = 4'b0000;
#5
A = 4'b1111;
B = 4'b0001;
#5
A = 4'b1111;
B = 4'b0010;
#5
A = 4'b1111;
B = 4'b0011;
#5
A = 4'b1111;
B = 4'b0100;
#5
A = 4'b1111;
B = 4'b0101;
#5
A = 4'b1111;
B = 4'b0110;
#5
A = 4'b1111;
B = 4'b0111;
#5
A = 4'b1111;
B = 4'b1000;
#5
A = 4'b1111;
B = 4'b1001;
#5
A = 4'b1111;
B = 4'b1010;
#5
A = 4'b1111;
B = 4'b1011;
#5
A = 4'b1111;
B = 4'b1100;
#5
A = 4'b1111;
B = 4'b1101;
#5
A = 4'b1111;
B = 4'b1110;
#5
A = 4'b1111;
B = 4'b1111;

end
endmodule

// iverilog -o run test.v
// vvp run
// gtkwave multiplier_tb.vcd