magic
tech scmos
timestamp 1669634335
<< metal1 >>
rect 54 1391 57 1417
<< metal2 >>
rect 135 1433 1009 1436
rect 58 1417 917 1420
rect 914 1275 917 1417
rect 1006 1275 1009 1433
<< polycontact >>
rect 54 1387 58 1391
<< m2contact >>
rect 54 1417 58 1421
use 4bit_multiplier  4bit_multiplier_0
timestamp 1669623720
transform 1 0 0 0 1 978
box 0 -978 1227 411
<< end >>
