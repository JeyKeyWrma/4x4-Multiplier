* SPICE3 file created from 4bit_adder.ext - technology: scmos

.option scale=1u

M1000 full_adder_1/Cin full_adder_0/or_0/inverter_0/input VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=40 pd=26 as=3040 ps=1976
M1001 full_adder_1/Cin full_adder_0/or_0/inverter_0/input GND Gnd nfet w=4 l=2
+  ad=20 pd=18 as=880 ps=792
M1002 full_adder_0/or_0/inverter_0/input full_adder_0/or_0/input2 full_adder_0/or_0/a_3_n6# full_adder_0/w_556_43# pfet w=8 l=2
+  ad=40 pd=26 as=80 ps=52
M1003 full_adder_0/or_0/a_3_n6# full_adder_0/or_0/input1 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 full_adder_0/or_0/inverter_0/input full_adder_0/or_0/input2 GND Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1005 full_adder_0/or_0/inverter_0/input full_adder_0/or_0/input1 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 full_adder_0/half_adder_1/nand_0/out full_adder_0/half_adder_1/input1 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1007 full_adder_0/half_adder_1/nand_0/out full_adder_0/half_adder_1/nand_2/input2 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 full_adder_0/half_adder_1/nand_0/out full_adder_0/half_adder_1/input1 full_adder_0/half_adder_1/nand_0/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1009 full_adder_0/half_adder_1/nand_0/a_3_n27# full_adder_0/half_adder_1/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 S1 full_adder_0/half_adder_1/nand_1/input2 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1011 S1 full_adder_0/half_adder_1/nand_0/out VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 S1 full_adder_0/half_adder_1/nand_1/input2 full_adder_0/half_adder_1/nand_1/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1013 full_adder_0/half_adder_1/nand_1/a_3_n27# full_adder_0/half_adder_1/nand_0/out GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 full_adder_0/or_0/input1 full_adder_0/half_adder_1/nand_2/input2 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1015 full_adder_0/or_0/input1 full_adder_0/half_adder_1/nand_2/input2 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 full_adder_0/or_0/input1 full_adder_0/half_adder_1/nand_2/input2 full_adder_0/half_adder_1/nand_2/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1017 full_adder_0/half_adder_1/nand_2/a_3_n27# full_adder_0/half_adder_1/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 full_adder_0/half_adder_1/nand_2/input2 full_adder_0/Cin VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1019 full_adder_0/half_adder_1/a_59_n27# full_adder_0/half_adder_1/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1020 full_adder_0/half_adder_1/nand_2/input2 full_adder_0/half_adder_1/input1 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1021 full_adder_0/half_adder_1/nand_1/input2 full_adder_0/Cin full_adder_0/half_adder_1/a_59_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1022 full_adder_0/half_adder_1/nand_2/input2 full_adder_0/Cin full_adder_0/half_adder_1/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1023 full_adder_0/half_adder_1/a_3_n27# full_adder_0/half_adder_1/input1 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 full_adder_0/half_adder_1/nand_1/input2 full_adder_0/half_adder_1/nand_2/input2 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1025 full_adder_0/half_adder_1/nand_1/input2 full_adder_0/Cin VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 full_adder_0/half_adder_0/nand_0/out A1 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1027 full_adder_0/half_adder_0/nand_0/out full_adder_0/half_adder_0/nand_2/input2 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 full_adder_0/half_adder_0/nand_0/out A1 full_adder_0/half_adder_0/nand_0/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1029 full_adder_0/half_adder_0/nand_0/a_3_n27# full_adder_0/half_adder_0/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 full_adder_0/half_adder_1/input1 full_adder_0/half_adder_0/nand_1/input2 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1031 full_adder_0/half_adder_1/input1 full_adder_0/half_adder_0/nand_0/out VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 full_adder_0/half_adder_1/input1 full_adder_0/half_adder_0/nand_1/input2 full_adder_0/half_adder_0/nand_1/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1033 full_adder_0/half_adder_0/nand_1/a_3_n27# full_adder_0/half_adder_0/nand_0/out GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 full_adder_0/or_0/input2 full_adder_0/half_adder_0/nand_2/input2 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1035 full_adder_0/or_0/input2 full_adder_0/half_adder_0/nand_2/input2 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 full_adder_0/or_0/input2 full_adder_0/half_adder_0/nand_2/input2 full_adder_0/half_adder_0/nand_2/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1037 full_adder_0/half_adder_0/nand_2/a_3_n27# full_adder_0/half_adder_0/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 full_adder_0/half_adder_0/nand_2/input2 B1 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1039 full_adder_0/half_adder_0/a_59_n27# full_adder_0/half_adder_0/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1040 full_adder_0/half_adder_0/nand_2/input2 A1 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 full_adder_0/half_adder_0/nand_1/input2 B1 full_adder_0/half_adder_0/a_59_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1042 full_adder_0/half_adder_0/nand_2/input2 B1 full_adder_0/half_adder_0/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1043 full_adder_0/half_adder_0/a_3_n27# A1 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 full_adder_0/half_adder_0/nand_1/input2 full_adder_0/half_adder_0/nand_2/input2 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1045 full_adder_0/half_adder_0/nand_1/input2 B1 VDD full_adder_0/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 full_adder_2/Cin full_adder_1/or_0/inverter_0/input VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1047 full_adder_2/Cin full_adder_1/or_0/inverter_0/input GND Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1048 full_adder_1/or_0/inverter_0/input full_adder_1/or_0/input2 full_adder_1/or_0/a_3_n6# full_adder_1/w_556_43# pfet w=8 l=2
+  ad=40 pd=26 as=80 ps=52
M1049 full_adder_1/or_0/a_3_n6# full_adder_1/or_0/input1 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 full_adder_1/or_0/inverter_0/input full_adder_1/or_0/input2 GND Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1051 full_adder_1/or_0/inverter_0/input full_adder_1/or_0/input1 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 full_adder_1/half_adder_1/nand_0/out full_adder_1/half_adder_1/input1 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1053 full_adder_1/half_adder_1/nand_0/out full_adder_1/half_adder_1/nand_2/input2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 full_adder_1/half_adder_1/nand_0/out full_adder_1/half_adder_1/input1 full_adder_1/half_adder_1/nand_0/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1055 full_adder_1/half_adder_1/nand_0/a_3_n27# full_adder_1/half_adder_1/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 S2 full_adder_1/half_adder_1/nand_1/input2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1057 S2 full_adder_1/half_adder_1/nand_0/out VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1058 S2 full_adder_1/half_adder_1/nand_1/input2 full_adder_1/half_adder_1/nand_1/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1059 full_adder_1/half_adder_1/nand_1/a_3_n27# full_adder_1/half_adder_1/nand_0/out GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 full_adder_1/or_0/input1 full_adder_1/half_adder_1/nand_2/input2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1061 full_adder_1/or_0/input1 full_adder_1/half_adder_1/nand_2/input2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 full_adder_1/or_0/input1 full_adder_1/half_adder_1/nand_2/input2 full_adder_1/half_adder_1/nand_2/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1063 full_adder_1/half_adder_1/nand_2/a_3_n27# full_adder_1/half_adder_1/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 full_adder_1/half_adder_1/nand_2/input2 full_adder_1/Cin VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1065 full_adder_1/half_adder_1/a_59_n27# full_adder_1/half_adder_1/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1066 full_adder_1/half_adder_1/nand_2/input2 full_adder_1/half_adder_1/input1 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 full_adder_1/half_adder_1/nand_1/input2 full_adder_1/Cin full_adder_1/half_adder_1/a_59_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1068 full_adder_1/half_adder_1/nand_2/input2 full_adder_1/Cin full_adder_1/half_adder_1/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1069 full_adder_1/half_adder_1/a_3_n27# full_adder_1/half_adder_1/input1 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 full_adder_1/half_adder_1/nand_1/input2 full_adder_1/half_adder_1/nand_2/input2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1071 full_adder_1/half_adder_1/nand_1/input2 full_adder_1/Cin VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1072 full_adder_1/half_adder_0/nand_0/out A2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1073 full_adder_1/half_adder_0/nand_0/out full_adder_1/half_adder_0/nand_2/input2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 full_adder_1/half_adder_0/nand_0/out A2 full_adder_1/half_adder_0/nand_0/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1075 full_adder_1/half_adder_0/nand_0/a_3_n27# full_adder_1/half_adder_0/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 full_adder_1/half_adder_1/input1 full_adder_1/half_adder_0/nand_1/input2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1077 full_adder_1/half_adder_1/input1 full_adder_1/half_adder_0/nand_0/out VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 full_adder_1/half_adder_1/input1 full_adder_1/half_adder_0/nand_1/input2 full_adder_1/half_adder_0/nand_1/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1079 full_adder_1/half_adder_0/nand_1/a_3_n27# full_adder_1/half_adder_0/nand_0/out GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1080 full_adder_1/or_0/input2 full_adder_1/half_adder_0/nand_2/input2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1081 full_adder_1/or_0/input2 full_adder_1/half_adder_0/nand_2/input2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 full_adder_1/or_0/input2 full_adder_1/half_adder_0/nand_2/input2 full_adder_1/half_adder_0/nand_2/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1083 full_adder_1/half_adder_0/nand_2/a_3_n27# full_adder_1/half_adder_0/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1084 full_adder_1/half_adder_0/nand_2/input2 B2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1085 full_adder_1/half_adder_0/a_59_n27# full_adder_1/half_adder_0/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1086 full_adder_1/half_adder_0/nand_2/input2 A2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 full_adder_1/half_adder_0/nand_1/input2 B2 full_adder_1/half_adder_0/a_59_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1088 full_adder_1/half_adder_0/nand_2/input2 B2 full_adder_1/half_adder_0/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1089 full_adder_1/half_adder_0/a_3_n27# A2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 full_adder_1/half_adder_0/nand_1/input2 full_adder_1/half_adder_0/nand_2/input2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1091 full_adder_1/half_adder_0/nand_1/input2 B2 VDD full_adder_1/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1092 C_OUT full_adder_2/or_0/inverter_0/input VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1093 C_OUT full_adder_2/or_0/inverter_0/input GND Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1094 full_adder_2/or_0/inverter_0/input full_adder_2/or_0/input2 full_adder_2/or_0/a_3_n6# full_adder_2/w_556_43# pfet w=8 l=2
+  ad=40 pd=26 as=80 ps=52
M1095 full_adder_2/or_0/a_3_n6# full_adder_2/or_0/input1 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 full_adder_2/or_0/inverter_0/input full_adder_2/or_0/input2 GND Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1097 full_adder_2/or_0/inverter_0/input full_adder_2/or_0/input1 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1098 full_adder_2/half_adder_1/nand_0/out full_adder_2/half_adder_1/input1 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1099 full_adder_2/half_adder_1/nand_0/out full_adder_2/half_adder_1/nand_2/input2 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 full_adder_2/half_adder_1/nand_0/out full_adder_2/half_adder_1/input1 full_adder_2/half_adder_1/nand_0/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1101 full_adder_2/half_adder_1/nand_0/a_3_n27# full_adder_2/half_adder_1/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 S3 full_adder_2/half_adder_1/nand_1/input2 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1103 S3 full_adder_2/half_adder_1/nand_0/out VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1104 S3 full_adder_2/half_adder_1/nand_1/input2 full_adder_2/half_adder_1/nand_1/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1105 full_adder_2/half_adder_1/nand_1/a_3_n27# full_adder_2/half_adder_1/nand_0/out GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1106 full_adder_2/or_0/input1 full_adder_2/half_adder_1/nand_2/input2 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1107 full_adder_2/or_0/input1 full_adder_2/half_adder_1/nand_2/input2 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1108 full_adder_2/or_0/input1 full_adder_2/half_adder_1/nand_2/input2 full_adder_2/half_adder_1/nand_2/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1109 full_adder_2/half_adder_1/nand_2/a_3_n27# full_adder_2/half_adder_1/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 full_adder_2/half_adder_1/nand_2/input2 full_adder_2/Cin VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1111 full_adder_2/half_adder_1/a_59_n27# full_adder_2/half_adder_1/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1112 full_adder_2/half_adder_1/nand_2/input2 full_adder_2/half_adder_1/input1 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 full_adder_2/half_adder_1/nand_1/input2 full_adder_2/Cin full_adder_2/half_adder_1/a_59_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1114 full_adder_2/half_adder_1/nand_2/input2 full_adder_2/Cin full_adder_2/half_adder_1/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1115 full_adder_2/half_adder_1/a_3_n27# full_adder_2/half_adder_1/input1 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 full_adder_2/half_adder_1/nand_1/input2 full_adder_2/half_adder_1/nand_2/input2 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1117 full_adder_2/half_adder_1/nand_1/input2 full_adder_2/Cin VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1118 full_adder_2/half_adder_0/nand_0/out A3 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1119 full_adder_2/half_adder_0/nand_0/out full_adder_2/half_adder_0/nand_2/input2 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 full_adder_2/half_adder_0/nand_0/out A3 full_adder_2/half_adder_0/nand_0/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1121 full_adder_2/half_adder_0/nand_0/a_3_n27# full_adder_2/half_adder_0/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 full_adder_2/half_adder_1/input1 full_adder_2/half_adder_0/nand_1/input2 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1123 full_adder_2/half_adder_1/input1 full_adder_2/half_adder_0/nand_0/out VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 full_adder_2/half_adder_1/input1 full_adder_2/half_adder_0/nand_1/input2 full_adder_2/half_adder_0/nand_1/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1125 full_adder_2/half_adder_0/nand_1/a_3_n27# full_adder_2/half_adder_0/nand_0/out GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1126 full_adder_2/or_0/input2 full_adder_2/half_adder_0/nand_2/input2 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1127 full_adder_2/or_0/input2 full_adder_2/half_adder_0/nand_2/input2 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 full_adder_2/or_0/input2 full_adder_2/half_adder_0/nand_2/input2 full_adder_2/half_adder_0/nand_2/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1129 full_adder_2/half_adder_0/nand_2/a_3_n27# full_adder_2/half_adder_0/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 full_adder_2/half_adder_0/nand_2/input2 B3 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1131 full_adder_2/half_adder_0/a_59_n27# full_adder_2/half_adder_0/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1132 full_adder_2/half_adder_0/nand_2/input2 A3 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1133 full_adder_2/half_adder_0/nand_1/input2 B3 full_adder_2/half_adder_0/a_59_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1134 full_adder_2/half_adder_0/nand_2/input2 B3 full_adder_2/half_adder_0/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1135 full_adder_2/half_adder_0/a_3_n27# A3 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 full_adder_2/half_adder_0/nand_1/input2 full_adder_2/half_adder_0/nand_2/input2 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1137 full_adder_2/half_adder_0/nand_1/input2 B3 VDD full_adder_2/w_556_43# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1138 half_adder_0/nand_0/out A0 VDD half_adder_0/w_n10_n12# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1139 half_adder_0/nand_0/out half_adder_0/nand_2/input2 VDD half_adder_0/w_n10_n12# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 half_adder_0/nand_0/out A0 half_adder_0/nand_0/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1141 half_adder_0/nand_0/a_3_n27# half_adder_0/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 S0 half_adder_0/nand_1/input2 VDD half_adder_0/w_n10_n12# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1143 S0 half_adder_0/nand_0/out VDD half_adder_0/w_n10_n12# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 S0 half_adder_0/nand_1/input2 half_adder_0/nand_1/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1145 half_adder_0/nand_1/a_3_n27# half_adder_0/nand_0/out GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 full_adder_0/Cin half_adder_0/nand_2/input2 VDD half_adder_0/w_n10_n12# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1147 full_adder_0/Cin half_adder_0/nand_2/input2 VDD half_adder_0/w_n10_n12# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 full_adder_0/Cin half_adder_0/nand_2/input2 half_adder_0/nand_2/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1149 half_adder_0/nand_2/a_3_n27# half_adder_0/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1150 half_adder_0/nand_2/input2 B0 VDD half_adder_0/w_n10_n12# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1151 half_adder_0/a_59_n27# half_adder_0/nand_2/input2 GND Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1152 half_adder_0/nand_2/input2 A0 VDD half_adder_0/w_n10_n12# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1153 half_adder_0/nand_1/input2 B0 half_adder_0/a_59_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1154 half_adder_0/nand_2/input2 B0 half_adder_0/a_3_n27# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1155 half_adder_0/a_3_n27# A0 GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1156 half_adder_0/nand_1/input2 half_adder_0/nand_2/input2 VDD half_adder_0/w_n10_n12# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1157 half_adder_0/nand_1/input2 B0 VDD half_adder_0/w_n10_n12# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
C0 full_adder_1/Cin full_adder_1/w_556_43# 6.35fF
C1 full_adder_0/w_556_43# full_adder_0/half_adder_0/nand_2/input2 14.96fF
C2 full_adder_0/w_556_43# full_adder_0/or_0/input1 5.43fF
C3 full_adder_1/half_adder_1/input1 full_adder_1/w_556_43# 13.37fF
C4 full_adder_2/w_556_43# full_adder_2/or_0/input1 5.43fF
C5 full_adder_2/w_556_43# full_adder_2/half_adder_1/nand_1/input2 5.43fF
C6 half_adder_0/w_n10_n12# B0 6.35fF
C7 half_adder_0/w_n10_n12# S0 2.26fF
C8 full_adder_0/w_556_43# VDD 24.82fF
C9 full_adder_0/w_556_43# full_adder_0/Cin 6.35fF
C10 full_adder_2/Cin full_adder_2/half_adder_1/input1 2.28fF
C11 full_adder_1/w_556_43# S2 2.26fF
C12 full_adder_0/w_556_43# B1 6.35fF
C13 half_adder_0/w_n10_n12# VDD 11.28fF
C14 full_adder_0/w_556_43# full_adder_0/or_0/inverter_0/input 4.30fF
C15 half_adder_0/w_n10_n12# full_adder_0/Cin 2.26fF
C16 full_adder_1/w_556_43# A2 6.35fF
C17 full_adder_2/w_556_43# B3 6.35fF
C18 full_adder_2/w_556_43# full_adder_2/half_adder_0/nand_0/out 5.43fF
C19 full_adder_0/w_556_43# full_adder_0/half_adder_1/input1 13.37fF
C20 full_adder_0/w_556_43# full_adder_0/half_adder_1/nand_1/input2 5.43fF
C21 full_adder_1/or_0/input1 full_adder_1/w_556_43# 5.43fF
C22 full_adder_2/w_556_43# VDD 24.82fF
C23 full_adder_1/w_556_43# full_adder_1/or_0/inverter_0/input 4.30fF
C24 full_adder_0/w_556_43# full_adder_0/or_0/a_3_n6# 6.39fF
C25 half_adder_0/w_n10_n12# half_adder_0/nand_0/out 5.43fF
C26 full_adder_2/w_556_43# full_adder_2/half_adder_1/nand_2/input2 14.96fF
C27 full_adder_1/half_adder_0/nand_0/out full_adder_1/w_556_43# 5.43fF
C28 full_adder_1/or_0/input2 full_adder_1/w_556_43# 5.43fF
C29 full_adder_1/w_556_43# full_adder_1/half_adder_1/nand_2/input2 14.96fF
C30 full_adder_2/w_556_43# full_adder_2/or_0/inverter_0/input 4.30fF
C31 full_adder_0/w_556_43# A1 6.35fF
C32 full_adder_1/half_adder_1/nand_1/input2 full_adder_1/w_556_43# 5.43fF
C33 full_adder_0/w_556_43# full_adder_0/half_adder_0/nand_1/input2 5.43fF
C34 full_adder_2/w_556_43# full_adder_2/half_adder_0/nand_1/input2 5.43fF
C35 full_adder_0/w_556_43# S1 2.26fF
C36 full_adder_2/w_556_43# full_adder_2/half_adder_1/nand_0/out 5.43fF
C37 half_adder_0/w_n10_n12# A0 6.35fF
C38 full_adder_2/w_556_43# full_adder_2/half_adder_0/nand_2/input2 14.96fF
C39 full_adder_2/w_556_43# full_adder_2/or_0/a_3_n6# 6.39fF
C40 full_adder_1/w_556_43# full_adder_1/half_adder_0/nand_1/input2 5.43fF
C41 full_adder_2/w_556_43# A3 6.35fF
C42 full_adder_1/half_adder_1/nand_0/out full_adder_1/w_556_43# 5.43fF
C43 full_adder_0/w_556_43# full_adder_0/half_adder_0/nand_0/out 5.43fF
C44 full_adder_2/w_556_43# full_adder_2/or_0/input2 5.43fF
C45 full_adder_0/w_556_43# full_adder_0/half_adder_1/nand_2/input2 14.96fF
C46 half_adder_0/nand_2/input2 half_adder_0/w_n10_n12# 14.96fF
C47 full_adder_2/w_556_43# full_adder_2/Cin 6.35fF
C48 VDD full_adder_1/w_556_43# 24.82fF
C49 full_adder_1/w_556_43# B2 6.35fF
C50 full_adder_0/w_556_43# full_adder_0/or_0/input2 5.43fF
C51 full_adder_1/or_0/a_3_n6# full_adder_1/w_556_43# 6.39fF
C52 half_adder_0/w_n10_n12# half_adder_0/nand_1/input2 5.43fF
C53 full_adder_2/w_556_43# S3 2.26fF
C54 full_adder_0/w_556_43# full_adder_0/half_adder_1/nand_0/out 5.43fF
C55 full_adder_2/w_556_43# full_adder_2/half_adder_1/input1 13.37fF
C56 full_adder_1/half_adder_0/nand_2/input2 full_adder_1/w_556_43# 14.96fF
C57 half_adder_0/a_59_n27# Gnd 3.20fF
C58 half_adder_0/a_3_n27# Gnd 3.20fF
C59 B0 Gnd 7.57fF
C60 half_adder_0/nand_2/a_3_n27# Gnd 3.20fF
C61 half_adder_0/nand_1/a_3_n27# Gnd 3.20fF
C62 S0 Gnd 7.99fF
C63 half_adder_0/nand_1/input2 Gnd 33.30fF
C64 half_adder_0/nand_0/out Gnd 18.47fF
C65 half_adder_0/nand_0/a_3_n27# Gnd 3.20fF
C66 A0 Gnd 57.53fF
C67 half_adder_0/nand_2/input2 Gnd 22.89fF
C68 full_adder_2/half_adder_0/a_59_n27# Gnd 3.20fF
C69 full_adder_2/half_adder_0/a_3_n27# Gnd 3.20fF
C70 B3 Gnd 8.60fF
C71 full_adder_2/half_adder_0/nand_2/a_3_n27# Gnd 3.20fF
C72 GND Gnd 529.27fF
C73 full_adder_2/or_0/input2 Gnd 31.72fF
C74 full_adder_2/half_adder_0/nand_1/a_3_n27# Gnd 3.20fF
C75 full_adder_2/half_adder_1/input1 Gnd 91.67fF
C76 full_adder_2/half_adder_0/nand_1/input2 Gnd 33.30fF
C77 full_adder_2/half_adder_0/nand_0/out Gnd 18.47fF
C78 full_adder_2/half_adder_0/nand_0/a_3_n27# Gnd 3.20fF
C79 A3 Gnd 58.80fF
C80 full_adder_2/half_adder_0/nand_2/input2 Gnd 22.89fF
C81 full_adder_2/half_adder_1/a_59_n27# Gnd 3.20fF
C82 full_adder_2/half_adder_1/a_3_n27# Gnd 3.20fF
C83 full_adder_2/half_adder_1/nand_2/a_3_n27# Gnd 3.20fF
C84 full_adder_2/or_0/input1 Gnd 18.80fF
C85 full_adder_2/half_adder_1/nand_1/a_3_n27# Gnd 3.20fF
C86 S3 Gnd 10.86fF
C87 VDD Gnd 535.42fF
C88 full_adder_2/half_adder_1/nand_1/input2 Gnd 33.30fF
C89 full_adder_2/half_adder_1/nand_0/out Gnd 18.47fF
C90 full_adder_2/half_adder_1/nand_0/a_3_n27# Gnd 3.20fF
C91 full_adder_2/half_adder_1/nand_2/input2 Gnd 22.89fF
C92 C_OUT Gnd 6.82fF
C93 full_adder_2/or_0/inverter_0/input Gnd 22.12fF
C94 full_adder_1/half_adder_0/a_59_n27# Gnd 3.20fF
C95 full_adder_1/half_adder_0/a_3_n27# Gnd 3.20fF
C96 B2 Gnd 8.60fF
C97 full_adder_1/half_adder_0/nand_2/a_3_n27# Gnd 3.20fF
C98 full_adder_1/or_0/input2 Gnd 31.72fF
C99 full_adder_1/half_adder_0/nand_1/a_3_n27# Gnd 3.20fF
C100 full_adder_1/half_adder_1/input1 Gnd 91.67fF
C101 full_adder_1/half_adder_0/nand_1/input2 Gnd 33.30fF
C102 full_adder_1/half_adder_0/nand_0/out Gnd 18.47fF
C103 full_adder_1/half_adder_0/nand_0/a_3_n27# Gnd 3.20fF
C104 A2 Gnd 58.80fF
C105 full_adder_1/half_adder_0/nand_2/input2 Gnd 22.89fF
C106 full_adder_1/half_adder_1/a_59_n27# Gnd 3.20fF
C107 full_adder_1/half_adder_1/a_3_n27# Gnd 3.20fF
C108 full_adder_1/half_adder_1/nand_2/a_3_n27# Gnd 3.20fF
C109 full_adder_1/or_0/input1 Gnd 18.80fF
C110 full_adder_1/half_adder_1/nand_1/a_3_n27# Gnd 3.20fF
C111 S2 Gnd 10.86fF
C112 full_adder_1/half_adder_1/nand_1/input2 Gnd 33.30fF
C113 full_adder_1/half_adder_1/nand_0/out Gnd 18.47fF
C114 full_adder_1/half_adder_1/nand_0/a_3_n27# Gnd 3.20fF
C115 full_adder_1/half_adder_1/nand_2/input2 Gnd 22.89fF
C116 full_adder_2/Cin Gnd 38.55fF
C117 full_adder_1/or_0/inverter_0/input Gnd 22.12fF
C118 full_adder_0/half_adder_0/a_59_n27# Gnd 3.20fF
C119 full_adder_0/half_adder_0/a_3_n27# Gnd 3.20fF
C120 B1 Gnd 8.60fF
C121 full_adder_0/half_adder_0/nand_2/a_3_n27# Gnd 3.20fF
C122 full_adder_0/or_0/input2 Gnd 31.72fF
C123 full_adder_0/half_adder_0/nand_1/a_3_n27# Gnd 3.20fF
C124 full_adder_0/half_adder_1/input1 Gnd 91.67fF
C125 full_adder_0/half_adder_0/nand_1/input2 Gnd 33.30fF
C126 full_adder_0/half_adder_0/nand_0/out Gnd 18.47fF
C127 full_adder_0/half_adder_0/nand_0/a_3_n27# Gnd 3.20fF
C128 A1 Gnd 58.80fF
C129 full_adder_0/half_adder_0/nand_2/input2 Gnd 22.89fF
C130 full_adder_0/half_adder_1/a_59_n27# Gnd 3.20fF
C131 full_adder_0/half_adder_1/a_3_n27# Gnd 3.20fF
C132 full_adder_0/Cin Gnd 20.18fF
C133 full_adder_0/half_adder_1/nand_2/a_3_n27# Gnd 3.20fF
C134 full_adder_0/or_0/input1 Gnd 18.80fF
C135 full_adder_0/half_adder_1/nand_1/a_3_n27# Gnd 3.20fF
C136 S1 Gnd 11.10fF
C137 full_adder_0/half_adder_1/nand_1/input2 Gnd 33.30fF
C138 full_adder_0/half_adder_1/nand_0/out Gnd 18.47fF
C139 full_adder_0/half_adder_1/nand_0/a_3_n27# Gnd 3.20fF
C140 full_adder_0/half_adder_1/nand_2/input2 Gnd 22.89fF
C141 full_adder_1/Cin Gnd 39.24fF
C142 full_adder_0/or_0/inverter_0/input Gnd 22.12fF
