.include 22nm_MGK.pm
.param SUPPLY = 1

vDD VDD GND 'SUPPLY'

va input1 0 pulse 0 SUPPLY 10ns 100ps 100ps 5ns 20ns

vb input2 0 pulse 0 SUPPLY 0ns 100ps 100ps 10ns 20ns

.option scale = 0.01u

M1000 nand_0/out input1 vdd w_n10_n12# pmos w=8 l=2
+  ad=80 pd=52 as=400 ps=260
M1001 nand_0/out nand_2/input2 vdd w_n10_n12# pmos w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 nand_0/out input1 nand_0/a_3_n27# Gnd nmos w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1003 nand_0/a_3_n27# nand_2/input2 gnd Gnd nmos w=4 l=2
+  ad=0 pd=0 as=100 ps=90
M1004 SUM_HA nand_1/input2 vdd w_n10_n12# pmos w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1005 SUM_HA nand_0/out vdd w_n10_n12# pmos w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 SUM_HA nand_1/input2 nand_1/a_3_n27# Gnd nmos w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1007 nand_1/a_3_n27# nand_0/out gnd Gnd nmos w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 CARRY_HA nand_2/input2 vdd w_n10_n12# pmos w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1009 CARRY_HA nand_2/input2 vdd w_n10_n12# pmos w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 CARRY_HA nand_2/input2 nand_2/a_3_n27# Gnd nmos w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1011 nand_2/a_3_n27# nand_2/input2 gnd Gnd nmos w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 nand_2/input2 input2 vdd w_n10_n12# pmos w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1013 a_59_n27# nand_2/input2 gnd Gnd nmos w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1014 nand_2/input2 input1 vdd w_n10_n12# pmos w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 nand_1/input2 input2 a_59_n27# Gnd nmos w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1016 nand_2/input2 input2 a_3_n27# Gnd nmos w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1017 a_3_n27# input1 gnd Gnd nmos w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 nand_1/input2 nand_2/input2 vdd w_n10_n12# pmos w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1019 nand_1/input2 input2 vdd w_n10_n12# pmos w=8 l=2
+  ad=0 pd=0 as=0 ps=0

.tran 0.1ns 100ns
.control
run

plot v( SUM_HA)+4 v(CARRY_HA)+6 v(input1)+2 v(input2) 

.endc