magic
tech scmos
timestamp 1669378488
<< nwell >>
rect -10 -12 65 8
<< polysilicon >>
rect 1 2 3 11
rect 30 2 32 11
rect 1 -23 3 -6
rect 30 -23 32 -6
rect 54 -17 70 -15
rect 1 -35 3 -27
rect 30 -35 32 -27
<< ndiffusion >>
rect 0 -27 1 -23
rect 3 -27 4 -23
rect 29 -27 30 -23
rect 32 -27 33 -23
<< pdiffusion >>
rect 0 -6 1 2
rect 3 -6 4 2
rect 29 -6 30 2
rect 32 -6 33 2
<< metal1 >>
rect -12 12 65 16
rect -4 2 0 12
rect 8 -6 25 2
rect 33 -14 37 -6
rect 4 -15 37 -14
rect 4 -18 50 -15
rect 4 -23 8 -18
rect 33 -19 50 -18
rect 71 -17 92 -13
rect 33 -23 37 -19
rect -4 -36 0 -27
rect 25 -36 29 -27
rect 53 -36 57 -33
rect -4 -40 57 -36
<< ntransistor >>
rect 1 -27 3 -23
rect 30 -27 32 -23
<< ptransistor >>
rect 1 -6 3 2
rect 30 -6 32 2
<< polycontact >>
rect 50 -19 54 -15
<< ndcontact >>
rect -4 -27 0 -23
rect 4 -27 8 -23
rect 25 -27 29 -23
rect 33 -27 37 -23
<< pdcontact >>
rect -4 -6 0 2
rect 4 -6 8 2
rect 25 -6 29 2
rect 33 -6 37 2
use inverter  inverter_0
timestamp 1669373674
transform 1 0 67 0 1 0
box -14 -36 20 16
<< labels >>
rlabel polysilicon 2 -13 2 -13 1 input1
rlabel metal1 13 -38 13 -38 1 gnd
rlabel polysilicon 31 -13 31 -13 1 input2
rlabel metal1 2 13 2 13 5 vdd
rlabel metal1 90 -15 90 -15 7 out
<< end >>
